/*
 *  Copyright (C) 2018  Siddharth J <www.siddharth.pro>
 *
 *  Permission to use, copy, modify, and/or distribute this software for any
 *  purpose with or without fee is hereby granted, provided that the above
 *  copyright notice and this permission notice appear in all copies.
 *
 *  THE SOFTWARE IS PROVIDED "AS IS" AND THE AUTHOR DISCLAIMS ALL WARRANTIES
 *  WITH REGARD TO THIS SOFTWARE INCLUDING ALL IMPLIED WARRANTIES OF
 *  MERCHANTABILITY AND FITNESS. IN NO EVENT SHALL THE AUTHOR BE LIABLE FOR
 *  ANY SPECIAL, DIRECT, INDIRECT, OR CONSEQUENTIAL DAMAGES OR ANY DAMAGES
 *  WHATSOEVER RESULTING FROM LOSS OF USE, DATA OR PROFITS, WHETHER IN AN
 *  ACTION OF CONTRACT, NEGLIGENCE OR OTHER TORTIOUS ACTION, ARISING OUT OF
 *  OR IN CONNECTION WITH THE USE OR PERFORMANCE OF THIS SOFTWARE.
 *
 */
`include "defines.v"

module proRISC (clk,reset,Mem_OUT_test);
  
  input clk;
  input reset;
  output [7:0] Mem_OUT_test;
  wire [7:0] Mem_IN; 
  wire [7:0] Mem_OUT; 
  wire [7:0] Mem_ADDR;
  wire write;
  
  processor processing_unit(clk,reset,Mem_IN,Mem_OUT,Mem_ADDR,write);
  memory memory_unit(clk,Mem_IN,Mem_OUT,Mem_ADDR,write);
  assign Mem_OUT_test=Mem_OUT;
  
endmodule
